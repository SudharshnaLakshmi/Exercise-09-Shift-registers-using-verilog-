library verilog;
use verilog.vl_types.all;
entity pipo_vlg_check_tst is
    port(
        PO              : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end pipo_vlg_check_tst;
