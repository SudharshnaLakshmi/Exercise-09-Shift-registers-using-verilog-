library verilog;
use verilog.vl_types.all;
entity piso_vlg_vec_tst is
end piso_vlg_vec_tst;
