library verilog;
use verilog.vl_types.all;
entity sipo_vlg_vec_tst is
end sipo_vlg_vec_tst;
