library verilog;
use verilog.vl_types.all;
entity pipo_vlg_vec_tst is
end pipo_vlg_vec_tst;
